// lms_ctr.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module lms_ctr (
		input  wire        clk_clk,                                 //                              clk.clk
		input  wire [31:0] exfifo_if_d_export,                      //                      exfifo_if_d.export
		output wire        exfifo_if_rd_export,                     //                     exfifo_if_rd.export
		input  wire        exfifo_if_rdempty_export,                //                exfifo_if_rdempty.export
		output wire [31:0] exfifo_of_d_export,                      //                      exfifo_of_d.export
		output wire        exfifo_of_wr_export,                     //                     exfifo_of_wr.export
		input  wire        exfifo_of_wrfull_export,                 //                 exfifo_of_wrfull.export
		output wire        exfifo_rst_export,                       //                       exfifo_rst.export
		output wire [7:0]  leds_external_connection_export,         //         leds_external_connection.export
		output wire [3:0]  lms_ctr_gpio_external_connection_export, // lms_ctr_gpio_external_connection.export
		inout  wire        scl_exp_export,                          //                          scl_exp.export
		inout  wire        sda_exp_export,                          //                          sda_exp.export
		input  wire        spi_1_adf_external_MISO,                 //               spi_1_adf_external.MISO
		output wire        spi_1_adf_external_MOSI,                 //                                 .MOSI
		output wire        spi_1_adf_external_SCLK,                 //                                 .SCLK
		output wire        spi_1_adf_external_SS_n,                 //                                 .SS_n
		input  wire        spi_1_dac_external_MISO,                 //               spi_1_dac_external.MISO
		output wire        spi_1_dac_external_MOSI,                 //                                 .MOSI
		output wire        spi_1_dac_external_SCLK,                 //                                 .SCLK
		output wire        spi_1_dac_external_SS_n,                 //                                 .SS_n
		input  wire        spi_lms_external_MISO,                   //                 spi_lms_external.MISO
		output wire        spi_lms_external_MOSI,                   //                                 .MOSI
		output wire        spi_lms_external_SCLK,                   //                                 .SCLK
		output wire [4:0]  spi_lms_external_SS_n,                   //                                 .SS_n
		input  wire [7:0]  switch_external_connection_export        //       switch_external_connection.export
	);

	wire         nios2_cpu_debug_reset_request_reset;                                         // nios2_cpu:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1]
	wire         nios2_cpu_custom_instruction_master_readra;                                  // nios2_cpu:D_ci_readra -> nios2_cpu_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_a;                                       // nios2_cpu:D_ci_a -> nios2_cpu_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_b;                                       // nios2_cpu:D_ci_b -> nios2_cpu_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_cpu_custom_instruction_master_c;                                       // nios2_cpu:D_ci_c -> nios2_cpu_custom_instruction_master_translator:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_readrb;                                  // nios2_cpu:D_ci_readrb -> nios2_cpu_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios2_cpu_custom_instruction_master_ipending;                                // nios2_cpu:W_ci_ipending -> nios2_cpu_custom_instruction_master_translator:ci_slave_ipending
	wire   [7:0] nios2_cpu_custom_instruction_master_n;                                       // nios2_cpu:D_ci_n -> nios2_cpu_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_result;                                  // nios2_cpu_custom_instruction_master_translator:ci_slave_result -> nios2_cpu:E_ci_result
	wire         nios2_cpu_custom_instruction_master_estatus;                                 // nios2_cpu:W_ci_estatus -> nios2_cpu_custom_instruction_master_translator:ci_slave_estatus
	wire  [31:0] nios2_cpu_custom_instruction_master_datab;                                   // nios2_cpu:E_ci_datab -> nios2_cpu_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_dataa;                                   // nios2_cpu:E_ci_dataa -> nios2_cpu_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_writerc;                                 // nios2_cpu:D_ci_writerc -> nios2_cpu_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_result;        // nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_cpu_custom_instruction_master_translator:comb_ci_master_result
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra;        // nios2_cpu_custom_instruction_master_translator:comb_ci_master_readra -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_a;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_a -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_b;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_b -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb;        // nios2_cpu_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_c;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_c -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus;       // nios2_cpu_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending;      // nios2_cpu_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab;         // nios2_cpu_custom_instruction_master_translator:comb_ci_master_datab -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa;         // nios2_cpu_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc;       // nios2_cpu_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_n;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_n -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result;         // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra;         // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab;          // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result; // nios_custom_instr_bitswap_0:result -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab;  // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_bitswap_0:datab
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_bitswap_0:dataa
	wire  [31:0] nios2_cpu_data_master_readdata;                                              // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                                           // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                                           // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [16:0] nios2_cpu_data_master_address;                                               // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                                            // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                                  // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_write;                                                 // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                                             // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                                       // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                                    // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [16:0] nios2_cpu_instruction_master_address;                                        // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                                           // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect;                   // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_chipselect -> Av_FIFO_Int_0:chipselect
	wire  [31:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata;                     // Av_FIFO_Int_0:readdata -> mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address;                      // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_address -> Av_FIFO_Int_0:address
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read;                         // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_read -> Av_FIFO_Int_0:read
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write;                        // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_write -> Av_FIFO_Int_0:write
	wire  [31:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata;                    // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_writedata -> Av_FIFO_Int_0:writedata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect;                 // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata;                   // i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest;                // i2c_opencores_0:wb_ack_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address;                    // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write;                      // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata;                  // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;                        // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;                     // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;                     // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;                         // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;                            // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;                      // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;                           // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;                       // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_oc_mem_s1_chipselect;                                      // mm_interconnect_0:oc_mem_s1_chipselect -> oc_mem:chipselect
	wire  [31:0] mm_interconnect_0_oc_mem_s1_readdata;                                        // oc_mem:readdata -> mm_interconnect_0:oc_mem_s1_readdata
	wire  [12:0] mm_interconnect_0_oc_mem_s1_address;                                         // mm_interconnect_0:oc_mem_s1_address -> oc_mem:address
	wire   [3:0] mm_interconnect_0_oc_mem_s1_byteenable;                                      // mm_interconnect_0:oc_mem_s1_byteenable -> oc_mem:byteenable
	wire         mm_interconnect_0_oc_mem_s1_write;                                           // mm_interconnect_0:oc_mem_s1_write -> oc_mem:write
	wire  [31:0] mm_interconnect_0_oc_mem_s1_writedata;                                       // mm_interconnect_0:oc_mem_s1_writedata -> oc_mem:writedata
	wire         mm_interconnect_0_oc_mem_s1_clken;                                           // mm_interconnect_0:oc_mem_s1_clken -> oc_mem:clken
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                                        // switch:readdata -> mm_interconnect_0:switch_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                                         // mm_interconnect_0:switch_s1_address -> switch:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                        // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                          // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                           // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                                             // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                         // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_lms_ctr_gpio_s1_chipselect;                                // mm_interconnect_0:lms_ctr_gpio_s1_chipselect -> lms_ctr_gpio:chipselect
	wire  [31:0] mm_interconnect_0_lms_ctr_gpio_s1_readdata;                                  // lms_ctr_gpio:readdata -> mm_interconnect_0:lms_ctr_gpio_s1_readdata
	wire   [2:0] mm_interconnect_0_lms_ctr_gpio_s1_address;                                   // mm_interconnect_0:lms_ctr_gpio_s1_address -> lms_ctr_gpio:address
	wire         mm_interconnect_0_lms_ctr_gpio_s1_write;                                     // mm_interconnect_0:lms_ctr_gpio_s1_write -> lms_ctr_gpio:write_n
	wire  [31:0] mm_interconnect_0_lms_ctr_gpio_s1_writedata;                                 // mm_interconnect_0:lms_ctr_gpio_s1_writedata -> lms_ctr_gpio:writedata
	wire         mm_interconnect_0_spi_lms_spi_control_port_chipselect;                       // mm_interconnect_0:spi_lms_spi_control_port_chipselect -> spi_lms:spi_select
	wire  [15:0] mm_interconnect_0_spi_lms_spi_control_port_readdata;                         // spi_lms:data_to_cpu -> mm_interconnect_0:spi_lms_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_lms_spi_control_port_address;                          // mm_interconnect_0:spi_lms_spi_control_port_address -> spi_lms:mem_addr
	wire         mm_interconnect_0_spi_lms_spi_control_port_read;                             // mm_interconnect_0:spi_lms_spi_control_port_read -> spi_lms:read_n
	wire         mm_interconnect_0_spi_lms_spi_control_port_write;                            // mm_interconnect_0:spi_lms_spi_control_port_write -> spi_lms:write_n
	wire  [15:0] mm_interconnect_0_spi_lms_spi_control_port_writedata;                        // mm_interconnect_0:spi_lms_spi_control_port_writedata -> spi_lms:data_from_cpu
	wire         mm_interconnect_0_spi_1_dac_spi_control_port_chipselect;                     // mm_interconnect_0:spi_1_DAC_spi_control_port_chipselect -> spi_1_DAC:spi_select
	wire  [15:0] mm_interconnect_0_spi_1_dac_spi_control_port_readdata;                       // spi_1_DAC:data_to_cpu -> mm_interconnect_0:spi_1_DAC_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_1_dac_spi_control_port_address;                        // mm_interconnect_0:spi_1_DAC_spi_control_port_address -> spi_1_DAC:mem_addr
	wire         mm_interconnect_0_spi_1_dac_spi_control_port_read;                           // mm_interconnect_0:spi_1_DAC_spi_control_port_read -> spi_1_DAC:read_n
	wire         mm_interconnect_0_spi_1_dac_spi_control_port_write;                          // mm_interconnect_0:spi_1_DAC_spi_control_port_write -> spi_1_DAC:write_n
	wire  [15:0] mm_interconnect_0_spi_1_dac_spi_control_port_writedata;                      // mm_interconnect_0:spi_1_DAC_spi_control_port_writedata -> spi_1_DAC:data_from_cpu
	wire         mm_interconnect_0_spi_1_adf_spi_control_port_chipselect;                     // mm_interconnect_0:spi_1_ADF_spi_control_port_chipselect -> spi_1_ADF:spi_select
	wire  [15:0] mm_interconnect_0_spi_1_adf_spi_control_port_readdata;                       // spi_1_ADF:data_to_cpu -> mm_interconnect_0:spi_1_ADF_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_1_adf_spi_control_port_address;                        // mm_interconnect_0:spi_1_ADF_spi_control_port_address -> spi_1_ADF:mem_addr
	wire         mm_interconnect_0_spi_1_adf_spi_control_port_read;                           // mm_interconnect_0:spi_1_ADF_spi_control_port_read -> spi_1_ADF:read_n
	wire         mm_interconnect_0_spi_1_adf_spi_control_port_write;                          // mm_interconnect_0:spi_1_ADF_spi_control_port_write -> spi_1_ADF:write_n
	wire  [15:0] mm_interconnect_0_spi_1_adf_spi_control_port_writedata;                      // mm_interconnect_0:spi_1_ADF_spi_control_port_writedata -> spi_1_ADF:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                                    // i2c_opencores_0:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                    // spi_lms:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                    // spi_1_DAC:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                    // spi_1_ADF:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_cpu_irq_irq;                                                           // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         rst_controller_reset_out_reset;                                              // rst_controller:reset_out -> [Av_FIFO_Int_0:rsi_nrst, i2c_opencores_0:wb_rst_i, irq_mapper:reset, leds:reset_n, lms_ctr_gpio:reset_n, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n, oc_mem:reset, rst_translator:in_reset, spi_1_ADF:reset_n, spi_1_DAC:reset_n, spi_lms:reset_n, switch:reset_n, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                          // rst_controller:reset_req -> [nios2_cpu:reset_req, oc_mem:reset_req, rst_translator:reset_req_in]

	avfifo #(
		.width (32)
	) av_fifo_int_0 (
		.clk            (clk_clk),                                                   //          clock.clk
		.address        (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect     (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect), //               .chipselect
		.write          (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write),      //               .write
		.writedata      (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata),  //               .writedata
		.read           (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read),       //               .read
		.readdata       (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata),   //               .readdata
		.rsi_nrst       (~rst_controller_reset_out_reset),                           //          reset.reset_n
		.coe_if_d       (exfifo_if_d_export),                                        //       cnd_if_d.export
		.coe_if_rd      (exfifo_if_rd_export),                                       //      cnd_if_rd.export
		.coe_of_wrfull  (exfifo_of_wrfull_export),                                   //  cnd_of_wrfull.export
		.coe_of_wr      (exfifo_of_wr_export),                                       //      cnd_of_wr.export
		.coe_of_d       (exfifo_of_d_export),                                        //       cnd_of_d.export
		.coe_if_rdempty (exfifo_if_rdempty_export),                                  // cnd_if_rdempty.export
		.coe_fifo_rst   (exfifo_rst_export)                                          //   cnd_fifo_rst.export
	);

	i2c_opencores i2c_opencores_0 (
		.wb_clk_i   (clk_clk),                                                      //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                               //      clock_reset.reset
		.scl_pad_io (scl_exp_export),                                               //       export_scl.export
		.sda_pad_io (sda_exp_export),                                               //       export_sda.export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                      // interrupt_sender.irq
	);

	lms_ctr_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_external_connection_export)       // external_connection.export
	);

	lms_ctr_lms_ctr_gpio lms_ctr_gpio (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_lms_ctr_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_lms_ctr_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_lms_ctr_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_lms_ctr_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_lms_ctr_gpio_s1_readdata),   //                    .readdata
		.out_port   (lms_ctr_gpio_external_connection_export)       // external_connection.export
	);

	lms_ctr_nios2_cpu nios2_cpu (
		.clk                                 (clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_result                         (nios2_cpu_custom_instruction_master_result),              // custom_instruction_master.result
		.D_ci_a                              (nios2_cpu_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (nios2_cpu_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (nios2_cpu_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (nios2_cpu_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (nios2_cpu_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (nios2_cpu_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (nios2_cpu_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (nios2_cpu_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (nios2_cpu_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (),                                                        //                          .clk
		.E_ci_multi_reset                    (),                                                        //                          .reset
		.E_ci_multi_reset_req                (),                                                        //                          .reset_req
		.W_ci_estatus                        (nios2_cpu_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (nios2_cpu_custom_instruction_master_ipending)             //                          .ipending
	);

	bitswap_qsys nios_custom_instr_bitswap_0 (
		.dataa  (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // s1.dataa
		.datab  (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //   .datab
		.result (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result)  //   .result
	);

	lms_ctr_oc_mem oc_mem (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_oc_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_oc_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_oc_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_oc_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_oc_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_oc_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_oc_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	lms_ctr_spi_1_ADF spi_1_adf (
		.clk           (clk_clk),                                                 //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                         //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_1_adf_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_1_adf_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_1_adf_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_1_adf_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_1_adf_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_1_adf_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                                //              irq.irq
		.MISO          (spi_1_adf_external_MISO),                                 //         external.export
		.MOSI          (spi_1_adf_external_MOSI),                                 //                 .export
		.SCLK          (spi_1_adf_external_SCLK),                                 //                 .export
		.SS_n          (spi_1_adf_external_SS_n)                                  //                 .export
	);

	lms_ctr_spi_1_DAC spi_1_dac (
		.clk           (clk_clk),                                                 //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                         //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_1_dac_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_1_dac_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_1_dac_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_1_dac_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_1_dac_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_1_dac_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                                //              irq.irq
		.MISO          (spi_1_dac_external_MISO),                                 //         external.export
		.MOSI          (spi_1_dac_external_MOSI),                                 //                 .export
		.SCLK          (spi_1_dac_external_SCLK),                                 //                 .export
		.SS_n          (spi_1_dac_external_SS_n)                                  //                 .export
	);

	lms_ctr_spi_lms spi_lms (
		.clk           (clk_clk),                                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_lms_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_lms_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_lms_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_lms_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_lms_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_lms_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver1_irq),                              //              irq.irq
		.MISO          (spi_lms_external_MISO),                                 //         external.export
		.MOSI          (spi_lms_external_MOSI),                                 //                 .export
		.SCLK          (spi_lms_external_SCLK),                                 //                 .export
		.SS_n          (spi_lms_external_SS_n)                                  //                 .export
	);

	lms_ctr_switch switch (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_s1_readdata), //                    .readdata
		.in_port  (switch_external_connection_export)     // external_connection.export
	);

	lms_ctr_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_cpu_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_cpu_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (nios2_cpu_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (nios2_cpu_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (nios2_cpu_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (nios2_cpu_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (nios2_cpu_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (nios2_cpu_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (nios2_cpu_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (nios2_cpu_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (nios2_cpu_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (nios2_cpu_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus          (nios2_cpu_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_done       (),                                                                       //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                   //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                   //    (terminated)
		.ci_slave_multi_result     (),                                                                       //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                            //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                   //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                               //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                               //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                               //    (terminated)
		.multi_ci_master_clk       (),                                                                       //    (terminated)
		.multi_ci_master_reset     (),                                                                       //    (terminated)
		.multi_ci_master_clken     (),                                                                       //    (terminated)
		.multi_ci_master_reset_req (),                                                                       //    (terminated)
		.multi_ci_master_start     (),                                                                       //    (terminated)
		.multi_ci_master_done      (1'b0),                                                                   //    (terminated)
		.multi_ci_master_dataa     (),                                                                       //    (terminated)
		.multi_ci_master_datab     (),                                                                       //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                                   //    (terminated)
		.multi_ci_master_n         (),                                                                       //    (terminated)
		.multi_ci_master_readra    (),                                                                       //    (terminated)
		.multi_ci_master_readrb    (),                                                                       //    (terminated)
		.multi_ci_master_writerc   (),                                                                       //    (terminated)
		.multi_ci_master_a         (),                                                                       //    (terminated)
		.multi_ci_master_b         (),                                                                       //    (terminated)
		.multi_ci_master_c         ()                                                                        //    (terminated)
	);

	lms_ctr_nios2_cpu_custom_instruction_master_comb_xconnect nios2_cpu_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (1)
	) nios2_cpu_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (),                                                                            // (terminated)
		.ci_master_readra    (),                                                                            // (terminated)
		.ci_master_readrb    (),                                                                            // (terminated)
		.ci_master_writerc   (),                                                                            // (terminated)
		.ci_master_a         (),                                                                            // (terminated)
		.ci_master_b         (),                                                                            // (terminated)
		.ci_master_c         (),                                                                            // (terminated)
		.ci_master_ipending  (),                                                                            // (terminated)
		.ci_master_estatus   (),                                                                            // (terminated)
		.ci_master_clk       (),                                                                            // (terminated)
		.ci_master_clken     (),                                                                            // (terminated)
		.ci_master_reset_req (),                                                                            // (terminated)
		.ci_master_reset     (),                                                                            // (terminated)
		.ci_master_start     (),                                                                            // (terminated)
		.ci_master_done      (1'b0),                                                                        // (terminated)
		.ci_slave_clk        (1'b0),                                                                        // (terminated)
		.ci_slave_clken      (1'b0),                                                                        // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                        // (terminated)
		.ci_slave_reset      (1'b0),                                                                        // (terminated)
		.ci_slave_start      (1'b0),                                                                        // (terminated)
		.ci_slave_done       ()                                                                             // (terminated)
	);

	lms_ctr_mm_interconnect_0 mm_interconnect_0 (
		.clk_main_clk_clk                            (clk_clk),                                                       //                          clk_main_clk.clk
		.nios2_cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // nios2_cpu_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address               (nios2_cpu_data_master_address),                                 //                 nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest           (nios2_cpu_data_master_waitrequest),                             //                                      .waitrequest
		.nios2_cpu_data_master_byteenable            (nios2_cpu_data_master_byteenable),                              //                                      .byteenable
		.nios2_cpu_data_master_read                  (nios2_cpu_data_master_read),                                    //                                      .read
		.nios2_cpu_data_master_readdata              (nios2_cpu_data_master_readdata),                                //                                      .readdata
		.nios2_cpu_data_master_write                 (nios2_cpu_data_master_write),                                   //                                      .write
		.nios2_cpu_data_master_writedata             (nios2_cpu_data_master_writedata),                               //                                      .writedata
		.nios2_cpu_data_master_debugaccess           (nios2_cpu_data_master_debugaccess),                             //                                      .debugaccess
		.nios2_cpu_instruction_master_address        (nios2_cpu_instruction_master_address),                          //          nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest    (nios2_cpu_instruction_master_waitrequest),                      //                                      .waitrequest
		.nios2_cpu_instruction_master_read           (nios2_cpu_instruction_master_read),                             //                                      .read
		.nios2_cpu_instruction_master_readdata       (nios2_cpu_instruction_master_readdata),                         //                                      .readdata
		.Av_FIFO_Int_0_avalon_slave_0_address        (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address),        //          Av_FIFO_Int_0_avalon_slave_0.address
		.Av_FIFO_Int_0_avalon_slave_0_write          (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write),          //                                      .write
		.Av_FIFO_Int_0_avalon_slave_0_read           (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read),           //                                      .read
		.Av_FIFO_Int_0_avalon_slave_0_readdata       (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata),       //                                      .readdata
		.Av_FIFO_Int_0_avalon_slave_0_writedata      (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata),      //                                      .writedata
		.Av_FIFO_Int_0_avalon_slave_0_chipselect     (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect),     //                                      .chipselect
		.i2c_opencores_0_avalon_slave_0_address      (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),      //        i2c_opencores_0_avalon_slave_0.address
		.i2c_opencores_0_avalon_slave_0_write        (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),        //                                      .write
		.i2c_opencores_0_avalon_slave_0_readdata     (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),     //                                      .readdata
		.i2c_opencores_0_avalon_slave_0_writedata    (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),    //                                      .writedata
		.i2c_opencores_0_avalon_slave_0_waitrequest  (~mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest), //                                      .waitrequest
		.i2c_opencores_0_avalon_slave_0_chipselect   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),   //                                      .chipselect
		.leds_s1_address                             (mm_interconnect_0_leds_s1_address),                             //                               leds_s1.address
		.leds_s1_write                               (mm_interconnect_0_leds_s1_write),                               //                                      .write
		.leds_s1_readdata                            (mm_interconnect_0_leds_s1_readdata),                            //                                      .readdata
		.leds_s1_writedata                           (mm_interconnect_0_leds_s1_writedata),                           //                                      .writedata
		.leds_s1_chipselect                          (mm_interconnect_0_leds_s1_chipselect),                          //                                      .chipselect
		.lms_ctr_gpio_s1_address                     (mm_interconnect_0_lms_ctr_gpio_s1_address),                     //                       lms_ctr_gpio_s1.address
		.lms_ctr_gpio_s1_write                       (mm_interconnect_0_lms_ctr_gpio_s1_write),                       //                                      .write
		.lms_ctr_gpio_s1_readdata                    (mm_interconnect_0_lms_ctr_gpio_s1_readdata),                    //                                      .readdata
		.lms_ctr_gpio_s1_writedata                   (mm_interconnect_0_lms_ctr_gpio_s1_writedata),                   //                                      .writedata
		.lms_ctr_gpio_s1_chipselect                  (mm_interconnect_0_lms_ctr_gpio_s1_chipselect),                  //                                      .chipselect
		.nios2_cpu_debug_mem_slave_address           (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),           //             nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write             (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),             //                                      .write
		.nios2_cpu_debug_mem_slave_read              (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),              //                                      .read
		.nios2_cpu_debug_mem_slave_readdata          (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),          //                                      .readdata
		.nios2_cpu_debug_mem_slave_writedata         (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),         //                                      .writedata
		.nios2_cpu_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),        //                                      .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest),       //                                      .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess),       //                                      .debugaccess
		.oc_mem_s1_address                           (mm_interconnect_0_oc_mem_s1_address),                           //                             oc_mem_s1.address
		.oc_mem_s1_write                             (mm_interconnect_0_oc_mem_s1_write),                             //                                      .write
		.oc_mem_s1_readdata                          (mm_interconnect_0_oc_mem_s1_readdata),                          //                                      .readdata
		.oc_mem_s1_writedata                         (mm_interconnect_0_oc_mem_s1_writedata),                         //                                      .writedata
		.oc_mem_s1_byteenable                        (mm_interconnect_0_oc_mem_s1_byteenable),                        //                                      .byteenable
		.oc_mem_s1_chipselect                        (mm_interconnect_0_oc_mem_s1_chipselect),                        //                                      .chipselect
		.oc_mem_s1_clken                             (mm_interconnect_0_oc_mem_s1_clken),                             //                                      .clken
		.spi_1_ADF_spi_control_port_address          (mm_interconnect_0_spi_1_adf_spi_control_port_address),          //            spi_1_ADF_spi_control_port.address
		.spi_1_ADF_spi_control_port_write            (mm_interconnect_0_spi_1_adf_spi_control_port_write),            //                                      .write
		.spi_1_ADF_spi_control_port_read             (mm_interconnect_0_spi_1_adf_spi_control_port_read),             //                                      .read
		.spi_1_ADF_spi_control_port_readdata         (mm_interconnect_0_spi_1_adf_spi_control_port_readdata),         //                                      .readdata
		.spi_1_ADF_spi_control_port_writedata        (mm_interconnect_0_spi_1_adf_spi_control_port_writedata),        //                                      .writedata
		.spi_1_ADF_spi_control_port_chipselect       (mm_interconnect_0_spi_1_adf_spi_control_port_chipselect),       //                                      .chipselect
		.spi_1_DAC_spi_control_port_address          (mm_interconnect_0_spi_1_dac_spi_control_port_address),          //            spi_1_DAC_spi_control_port.address
		.spi_1_DAC_spi_control_port_write            (mm_interconnect_0_spi_1_dac_spi_control_port_write),            //                                      .write
		.spi_1_DAC_spi_control_port_read             (mm_interconnect_0_spi_1_dac_spi_control_port_read),             //                                      .read
		.spi_1_DAC_spi_control_port_readdata         (mm_interconnect_0_spi_1_dac_spi_control_port_readdata),         //                                      .readdata
		.spi_1_DAC_spi_control_port_writedata        (mm_interconnect_0_spi_1_dac_spi_control_port_writedata),        //                                      .writedata
		.spi_1_DAC_spi_control_port_chipselect       (mm_interconnect_0_spi_1_dac_spi_control_port_chipselect),       //                                      .chipselect
		.spi_lms_spi_control_port_address            (mm_interconnect_0_spi_lms_spi_control_port_address),            //              spi_lms_spi_control_port.address
		.spi_lms_spi_control_port_write              (mm_interconnect_0_spi_lms_spi_control_port_write),              //                                      .write
		.spi_lms_spi_control_port_read               (mm_interconnect_0_spi_lms_spi_control_port_read),               //                                      .read
		.spi_lms_spi_control_port_readdata           (mm_interconnect_0_spi_lms_spi_control_port_readdata),           //                                      .readdata
		.spi_lms_spi_control_port_writedata          (mm_interconnect_0_spi_lms_spi_control_port_writedata),          //                                      .writedata
		.spi_lms_spi_control_port_chipselect         (mm_interconnect_0_spi_lms_spi_control_port_chipselect),         //                                      .chipselect
		.switch_s1_address                           (mm_interconnect_0_switch_s1_address),                           //                             switch_s1.address
		.switch_s1_readdata                          (mm_interconnect_0_switch_s1_readdata),                          //                                      .readdata
		.sysid_qsys_0_control_slave_address          (mm_interconnect_0_sysid_qsys_0_control_slave_address),          //            sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata         (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)          //                                      .readdata
	);

	lms_ctr_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_cpu_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_cpu_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
